`ifndef __utility_vh__
`define __utility_vh__

`define N 32
`define M 4

`endif